// Code your design here
module four_bit_pc(A_in, B_in, A, B, C, clk, Addr, SF, ZF,HLT, IP, OUTPORT, BYTE, SP);
  input [3:0]A_in;
  input [3:0]B_in;
  input [3:0]BYTE;
  input clk;
  
  
  reg carry = 0;
  reg [3:0]MEM[15:0];
  reg[3:0]STACK[15:0];
  reg load = 1;
  
  
  output reg [3:0]IP = 0;
  output reg [3:0]SP = 0;
  output reg[3:0]A, B, C, OUTPORT;
  output reg[3:0]Addr  = 0;
  output reg SF = 0;
  output reg ZF = 0;
  output reg HLT = 0;
  
  
  
  
  always @(posedge clk)
    begin
      MEM[0] 	= 4'b0100;
      MEM[1] 	= 4'b0110;
      MEM[2] 	= 4'b0100;
      MEM[3]	= 4'b0000;
      MEM[4] 	= 4'b0000;
      MEM[5] 	= 4'b0000;
      MEM[6] 	= 4'b1000;
      MEM[7] 	= 4'b0000;
      MEM[8] 	= 4'b0000;
      MEM[9] 	= 4'b0010;
      MEM[10] 	= 4'b1100;
      MEM[11] 	= 4'b0000;
      MEM[12] 	= 4'b0000;
      MEM[13] 	= 4'b1100;
      MEM[14] 	= 4'b0011;
      MEM[15] 	= 4'b1110;
		
		
		
		STACK[0] 	= 4'b0101;
		STACK[1] 	= 4'b0100;
		STACK[2] 	= 4'b0001;
		STACK[3] 	= 4'b0001;
		STACK[4] 	= 4'b0111;
		STACK[5] 	= 4'b0111;
		STACK[6] 	= 4'b0101;
		STACK[7] 	= 4'b0101;
		STACK[8] 	= 4'b0101;
		STACK[9] 	= 4'b0000;
		STACK[10] 	= 4'b0101;
		STACK[11] 	= 4'b0101;
		STACK[12] 	= 4'b0000;
		STACK[13] 	= 4'b0101;
		STACK[14] 	= 4'b0100;
		STACK[15] 	= 4'b0101;
		
      
		if (load == 1)
	     begin
		    A = A_in;
		    B = B_in;
		    load = 0;
		  end
		  
///////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////// Add A, B ////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////
      
      if (IP == 0)			
        begin
          {carry, C} = A + B; 
          A = C;
          C = 0;
          ZF = (A == 0)? 1:0;
          SF = (A < 0)? 1:0;
          
          IP = 1;
        end
		  
///////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////// Sub A, B ////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////
      else if (IP == 1)		
        begin
          {carry, C} = A - B; 
          A = C;
          C = 0;
          ZF = (A == 0)? 1:0;
          SF = (A < 0)? 1:0;
          
          IP = 2;
        end

		  
///////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////// XCHG B, A /////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////
      
      else if (IP == 2)		
        begin
          C = A;
          A = B;
          B = C;
          C = 0;
          
          ZF = (A == 0)?1:0;
          SF = (A < 0)?1:0;
          
          IP = 3;
        end
		  
////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////// mov B, [address] /////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////		  
      
      else if (IP == 3)		
         begin
           B = MEM[Addr];
           
           IP = 4;
         end

			
////////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////// out B ///////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////			
      else if (IP == 4)		
        begin
          OUTPORT = B;
          
          IP = 5;
        end
 
////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////// jnz Address ///////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////////////// 
      else if (IP == 5)		      
        begin
          if (ZF != 0)
            begin
              Addr = 8;
              IP = Addr;
            end
          else
            IP = 6;
        end

////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////  RCR A //////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////
		  
      else if (IP == 6)		 			
        begin
          C = (A>>1)+carry*8;			
			 A = C;
          
          IP = 7;
        end

////////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////// mov B, BYTE/////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////		  
      else if (IP == 7)		
        begin
          B = BYTE;
          
          IP = 8;
        end
////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////jmp Address //////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////


      else if (IP == 8)		
        begin
          Addr = 9;
          IP = Addr;
        end

////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////// push A ///////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////		  
      else if (IP == 9)		
        begin
          STACK[SP] = A;
          SP = SP + 1;
          ZF = (A == 0)?1:0;
          SF = (A<0) ? 1:0;
          
          IP = 10;
        end
      
////////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////// pop A	///////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////

      else if (IP == 10)		
        begin
          SP = SP - 1;
          A = STACK[SP];
          ZF = (STACK[SP] == 0)? 1:0;
          SF = (STACK[SP] < 0)? 1:0;
          
          IP = 11;
        end

////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////// CALL Addr/////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////
		  
      else if(IP == 11)		
        begin
          Addr = 13;
          STACK[SP] = IP;
          IP = Addr;
          SP = SP + 1;
        end

////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////// RET //////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////

      else if(IP == 12)		
        begin
          SP = SP - 1;
          IP = STACK[SP];
        end
		  
////////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////// xor A, [Addr] //////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////		  
      
      else if (IP == 13)		
        begin
          C = A^MEM[Addr];
          A = C;
          C = 0;
          ZF = (A == 0)?1:0;
          SF = (A<0)?1:0;
          
          IP = 14;
        end

///////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////test B, BYTE//////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////
		  
      else if (IP == 14)		
        begin
          C = B & BYTE;
          ZF = (C == 0)?1:0;
          SF = (C < 0)?1:0;
          C = 0;
          
          IP = 15;
        end
///////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////// HLT ///////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////      
      else if (IP == 15)		
        begin
          HLT = 1;
        end
            
      
      
      
    end
  
  
endmodule